/*******************************************************************************
 *
 * Copyright(C) 2008-2017 ERC CISST, Johns Hopkins University.
 *
 * This module measures the encoder pulse period by counting the edges of a
 * fixed fast clock (~3 MHz) between encoder pulses.  Each new encoder pulse
 * latches the current count and starts a new one.  From this measurement the
 * encoder period can be obtained by multiplying the number of counts by the
 * period of the fixed fast clock.
 *
 * Assumes counter will overflow if encoder moves too slowly.
 *
 * Revision history
 *     07/20/08    Paul Thienphrapa    Initial revision
 *     11/21/11    Paul Thienphrapa    Fix to use ticks+ as clock
 *     02/27/12    Paul Thienphrapa    Only count up due to unknown problem
 *     02/29/12    Zihan Chen          Fix implementation and debug module
 *     03/17/14    Peter Kazanzides    Update data every tick (dP = 4)
 *     04/07/17    Jie Ying Wu         Return only larger of cnter or cnter_latch
 */

module EncPeriod(
   input wire clk_fast,      // count this clock between encoder ticks
   input wire reset,         // global reset signal
   input wire ticks,         // encoder transition signal
   input wire dir,           // direction of the ticks
   output wire ticks_en,     // edge signal
   output reg[21:0] latched, // latched counter from last encoder event
   output reg[21:0] count,   // number clk_fast periods per tick
   output reg dir_changed,
   output reg overflowed
);

    // overflow value for unsigned 22-bit number
    parameter overflow = 22'h3FFFFF;


//------------------------------------------------------------------------------
// hardware description
//

// convert ticks to pulse
reg dir_r;      // dir start 
wire dir_diff;  // non-latched indication for direction change
reg ticks_r;    // previous ticks
assign ticks_en = ticks & (~ticks_r);
assign dir_diff = dir ^ dir_r;

always @(posedge clk_fast)
begin
   ticks_r <= ticks;
   dir_r <= dir;
end

// latch counter value
always @(posedge ticks_en or negedge reset)
begin
    if (reset == 0) begin
        latched <= 22'd0;
    end
    else begin
        latched <= count;
    end
end

// free-running counter 
always @(posedge clk_fast or posedge ticks_en or negedge reset) 
begin
   if (reset == 0 || ticks_en) begin
      count <= 22'd0;
      dir_changed <= 0;
      overflowed <= 0;
   end
   else if (dir_diff) begin
      dir_changed <= 1'b1;
   end
   else if (count != overflow) begin
      count <= count + 22'b1;
   end 
   else if (count == (overflow-22'b1)) begin
      overflowed <= 1'b0;
   end
end

endmodule


// ------------------------------------------------
// Quad Ticks Version 
// ------------------------------------------------
module EncPeriodQuad(
    input wire clk,           // sysclk
    input wire clk_fast,      // count this clock between encoder ticks
    input wire reset,         // global reset signal
    input wire a,             // quad encoder line a
    input wire b,             // quad encoder line b
    input wire dir,           // dir from EncQuad
    output reg[31:0] period,  // num of fast clock ticks
    output wire[31:0] acc      // [31:16] time since last edge, [15:0] estimated acc
);

    reg[1:0] mux;
    wire a_up_tick;
    wire a_dn_tick;
    wire b_up_tick;
    wire b_dn_tick;
    wire[21:0] a_up_latched;   // channel a up latched value
    wire[21:0] a_dn_latched;   // channel a dn latched value
    wire[21:0] b_up_latched;   // channel b up latched value
    wire[21:0] b_dn_latched;   // channel b dn latched value
    wire[21:0] a_up_counter;   // channel a up free running counter
    wire[21:0] a_dn_counter;   // channel a dn free running counter
    wire[21:0] b_up_counter;   // channel b up free running counter
    wire[21:0] b_dn_counter;   // channel b dn free running counter
    wire a_up_dir_changed;
    wire a_dn_dir_changed;
    wire b_up_dir_changed;
    wire b_dn_dir_changed;
    wire a_up_overflow;
    wire a_dn_overflow;
    wire b_up_overflow;
    wire b_dn_overflow;
    
//------------------------------------------------------------------------------
// hardware description
//

EncPeriod EncPerUpA(clk_fast, reset,  a, dir, a_up_tick, a_up_latched, a_up_counter, a_up_dir_changed, a_up_overflow);
EncPeriod EncPerDnA(clk_fast, reset, ~a, dir, a_dn_tick, a_dn_latched, a_dn_counter, a_dn_dir_changed, a_dn_overflow);
EncPeriod EncPerUpB(clk_fast, reset,  b, dir, b_up_tick, b_up_latched, b_up_counter, b_up_dir_changed, b_up_overflow);
EncPeriod EncPerDnB(clk_fast, reset, ~b, dir, b_dn_tick, b_dn_latched, b_dn_counter, b_dn_dir_changed, b_dn_overflow);

localparam[1:0] a_up = 2'b00;
localparam[1:0] a_dn = 2'b01;
localparam[1:0] b_up = 2'b10;
localparam[1:0] b_dn = 2'b11;

//Keep track of last 2 periods for acceleration and counter since last tick
reg[15:0] counter [1:6];

wire any_tick;
assign any_tick = a_up_tick | a_dn_tick | b_up_tick | b_dn_tick;

// Determine which edge is the most recent
always @(posedge any_tick)
begin
    if (a_up_tick) begin
        mux <= a_up;
    end
    else if (b_up_tick) begin
        mux <= b_up;    
    end    
    else if (a_dn_tick) begin
        mux <= a_dn;
    end
    else if (b_dn_tick) begin
        mux <= b_dn;
    end
    
end

always @(posedge clk_fast) begin
    if (any_tick) begin
        counter[1] <= 16'b0;
        counter[2] <= counter[1];
        counter[3] <= counter[2];
        counter[4] <= counter[3];
        counter[5] <= counter[4];
        counter[6] <= counter[5];
    end else if (counter[1] != 16'hFFFF) begin
        counter[1] <= counter[1] + 16'b1;
    end
end

assign acc[15:0] = counter[6];
assign acc[31:16] = counter[2]; 

// The following code returns the larger of (1) the most recent latched value (determined by mux)
// or (2) the free-running counter for the next expected encoder transition, based on direction, dir.
// Note that a direction change sets the free-running counter to overflow, so that will take priority
// over the latched value, which is reasonable behavior (i.e., a recent direction change should result
// in an estimated velocity of 0).
// From EncQuad.v:
//   dir 0 is A leading B  (cycle is Aup -> Bup -> Adown -> Bdown)
//   dir 1 is B leading A  (cycle is Bup -> Aup -> Bdown -> Adown)
always @(posedge clk_fast or negedge reset) begin
   if (reset == 0) begin
      period <= 32'd0;
   end
   
   else if (mux == a_up) begin  // A up
         period <= {1'b1, dir, a_up_dir_changed, a_up, a_up_overflow, 4'd0, a_up_latched};
   end

   else if (mux == b_up) begin  // B up
         period <= {1'b1, dir, b_up_dir_changed, b_up, b_up_overflow, 4'd0, b_up_latched};
   end

   else if (mux == a_dn) begin  // A down
         period <= {1'b1, dir, a_dn_dir_changed, a_dn, a_dn_overflow, 4'd0, a_dn_latched};
   end

   else if (mux == b_dn) begin  // B down
         period <= {1'b1, dir, b_dn_dir_changed, b_dn, b_dn_overflow, 4'd0, b_dn_latched};
   end
   
end

endmodule
